`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/18/2020 09:29:38 PM
// Design Name: 
// Module Name: HW_2_Nagelvoort_Ethan_Prob1_2always
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module HW_2_Nagelvoort_Ethan_Prob1_2always(

    );
endmodule
